////////////////////////////////////////////////////////////////////////////////
// Filename    : decoder_4to16.v
// Description : 
//
// Author      : Phu Vuong
// History     : Aug 15, 2023 : Initial     
//
////////////////////////////////////////////////////////////////////////////////
module decoder_4to16(
    //-----------------------
    //input
    en_i,
    in_i,
    //-----------------------
    //output
    out_o
);
    ////////////////////////////////////////////////////////////////////////////
    //param declaration
    ////////////////////////////////////////////////////////////////////////////
	
	
    ////////////////////////////////////////////////////////////////////////////
    //pin - port declaration
    ////////////////////////////////////////////////////////////////////////////
    input                               en_i;
    input   [3:0]                       in_i;
    output  [15:0]                      out_o;
    
    ////////////////////////////////////////////////////////////////////////////
    //wire - reg name declaration
    ////////////////////////////////////////////////////////////////////////////
    wire    [3:0]                       int_en;

    ////////////////////////////////////////////////////////////////////////////
    //design description
    ////////////////////////////////////////////////////////////////////////////
    decoder_2to4 decoder_2to4_ctrl(
        .en_i(en_i),
        .in_i(in_i[3:2]),
        .out_o(int_en[3:0])
    );

    decoder_2to4 decoder_2to4_00(
        .en_i(int_en[0]),
        .in_i(in_i[1:0]),
        .out_o(out_o[3:0])
    );

    decoder_2to4 decoder_2to4_01(
        .en_i(int_en[1]),
        .in_i(in_i[1:0]),
        .out_o(out_o[7:4])
    );

    decoder_2to4 decoder_2to4_02(
        .en_i(int_en[2]),
        .in_i(in_i[1:0]),
        .out_o(out_o[11:8])
    );

    decoder_2to4 decoder_2to4_03(
        .en_i(int_en[3]),
        .in_i(in_i[1:0]),
        .out_o(out_o[15:12])
    );
endmodule
