////////////////////////////////////////////////////////////////////////////////
// Filename    : decoder_2to4.v
// Description : 
//
// Author      : Phu Vuong
// History     : Aug 15, 2023 : Initial     
//
////////////////////////////////////////////////////////////////////////////////
module decoder_2to4(
    //-----------------------
    //input
    en_i,
    in_i,
    //-----------------------
    //output
    out_o
);
    ////////////////////////////////////////////////////////////////////////////
    //param declaration
    ////////////////////////////////////////////////////////////////////////////
	
	
    ////////////////////////////////////////////////////////////////////////////
    //pin - port declaration
    ////////////////////////////////////////////////////////////////////////////
    input                               en_i;
    input   [1:0]                       in_i;
    output  [3:0]                       out_o;
    
    ////////////////////////////////////////////////////////////////////////////
    //wire - reg name declaration
    ////////////////////////////////////////////////////////////////////////////


    ////////////////////////////////////////////////////////////////////////////
    //design description
    ////////////////////////////////////////////////////////////////////////////
    assign out_o[3] = en_i & in_i[1] & in_i[0];
    assign out_o[2] = en_i & in_i[1] & (~in_i[0]);
    assign out_o[1] = en_i & (~in_i[1]) & in_i[0];
    assign out_o[0] = en_i & (~in_i[1]) & (~in_i[0]);
endmodule
